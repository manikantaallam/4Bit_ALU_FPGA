library ieee;
use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;


entity ROM_Decimal_Equivalents is
  port (
        --clk     :in std_logic;
       -- reset   :in std_logic;

        --Address for ROM Data
        Cur_D_Val_Out :in integer range 0 to 255;
        

        --Output for Seven Segments // Shall portmap accordingly to the SSHandler component
        Cur_D_Val_SS_out :out std_logic_vector(23 downto 0)  --dp,g,f,e,d,c,b,a --dp,g,f,e,d,c,b,a --dp,g,f,e,d,c,b,a
         
  );
end ROM_Decimal_Equivalents;

architecture struct of ROM_Decimal_Equivalents is  


  type ROM is Array (0 to 255) of std_logic_vector(23 downto 0);  
  signal ROM_Data :ROM := (

    "110000001111111111111111" ,   --0 
    "111110011111111111111111" ,   --1 
    "101001001111111111111111" ,   --2 
    "101100001111111111111111" ,   --3 
    "100110011111111111111111" ,   --4 
    "100100101111111111111111" ,   --5 
    "100000101111111111111111" ,   --6 
    "111110001111111111111111" ,   --7 
    "100000001111111111111111" ,   --8 
    "100100001111111111111111" ,   --9 
    "110000001111100111111111" ,   --10 
    "111110011111100111111111" ,   --11 
    "101001001111100111111111" ,   --12 
    "101100001111100111111111" ,   --13 
    "100110011111100111111111" ,   --14 
    "100100101111100111111111" ,   --15 
    "100000101111100111111111" ,   --16 
    "111110001111100111111111" ,   --17 
    "100000001111100111111111" ,   --18 
    "100100001111100111111111" ,   --19 
    "110000001010010011111111" ,   --20 
    "111110011010010011111111" ,   --21 
    "101001001010010011111111" ,   --22 
    "101100001010010011111111" ,   --23 
    "100110011010010011111111" ,   --24 
    "100100101010010011111111" ,   --25 
    "100000101010010011111111" ,   --26 
    "111110001010010011111111" ,   --27 
    "100000001010010011111111" ,   --28 
    "100100001010010011111111" ,   --29 
    "110000001011000011111111" ,   --30 
    "111110011011000011111111" ,   --31 
    "101001001011000011111111" ,   --32 
    "101100001011000011111111" ,   --33 
    "100110011011000011111111" ,   --34 
    "100100101011000011111111" ,   --35 
    "100000101011000011111111" ,   --36 
    "111110001011000011111111" ,   --37 
    "100000001011000011111111" ,   --38 
    "100100001011000011111111" ,   --39 
    "110000001001100111111111" ,   --40 
    "111110011001100111111111" ,   --41 
    "101001001001100111111111" ,   --42 
    "101100001001100111111111" ,   --43 
    "100110011001100111111111" ,   --44 
    "100100101001100111111111" ,   --45 
    "100000101001100111111111" ,   --46 
    "111110001001100111111111" ,   --47 
    "100000001001100111111111" ,   --48 
    "100100001001100111111111" ,   --49 
    "110000001001001011111111" ,   --50 
    "111110011001001011111111" ,   --51 
    "101001001001001011111111" ,   --52 
    "101100001001001011111111" ,   --53 
    "100110011001001011111111" ,   --54 
    "100100101001001011111111" ,   --55 
    "100000101001001011111111" ,   --56 
    "111110001001001011111111" ,   --57 
    "100000001001001011111111" ,   --58 
    "100100001001001011111111" ,   --59 
    "110000001000001011111111" ,   --60 
    "111110011000001011111111" ,   --61 
    "101001001000001011111111" ,   --62 
    "101100001000001011111111" ,   --63 
    "100110011000001011111111" ,   --64 
    "100100101000001011111111" ,   --65 
    "100000101000001011111111" ,   --66 
    "111110001000001011111111" ,   --67 
    "100000001000001011111111" ,   --68 
    "100100001000001011111111" ,   --69 
    "110000001111100011111111" ,   --70 
    "111110011111100011111111" ,   --71 
    "101001001111100011111111" ,   --72 
    "101100001111100011111111" ,   --73 
    "100110011111100011111111" ,   --74 
    "100100101111100011111111" ,   --75 
    "100000101111100011111111" ,   --76 
    "111110001111100011111111" ,   --77 
    "100000001111100011111111" ,   --78 
    "100100001111100011111111" ,   --79 
    "110000001000000011111111" ,   --80 
    "111110011000000011111111" ,   --81 
    "101001001000000011111111" ,   --82 
    "101100001000000011111111" ,   --83 
    "100110011000000011111111" ,   --84 
    "100100101000000011111111" ,   --85 
    "100000101000000011111111" ,   --86 
    "111110001000000011111111" ,   --87 
    "100000001000000011111111" ,   --88 
    "100100001000000011111111" ,   --89 
    "110000001001000011111111" ,   --90 
    "111110011001000011111111" ,   --91 
    "101001001001000011111111" ,   --92 
    "101100001001000011111111" ,   --93 
    "100110011001000011111111" ,   --94 
    "100100101001000011111111" ,   --95 
    "100000101001000011111111" ,   --96 
    "111110001001000011111111" ,   --97 
    "100000001001000011111111" ,   --98 
    "100100001001000011111111" ,   --99 
    "110000001100000011111001" ,   --100 
    "111110011100000011111001" ,   --101 
    "101001001100000011111001" ,   --102 
    "101100001100000011111001" ,   --103 
    "100110011100000011111001" ,   --104 
    "100100101100000011111001" ,   --105 
    "100000101100000011111001" ,   --106 
    "111110001100000011111001" ,   --107 
    "100000001100000011111001" ,   --108 
    "100100001100000011111001" ,   --109 
    "110000001111100111111001" ,   --110 
    "111110011111100111111001" ,   --111 
    "101001001111100111111001" ,   --112 
    "101100001111100111111001" ,   --113 
    "100110011111100111111001" ,   --114 
    "100100101111100111111001" ,   --115 
    "100000101111100111111001" ,   --116 
    "111110001111100111111001" ,   --117 
    "100000001111100111111001" ,   --118 
    "100100001111100111111001" ,   --119 
    "110000001010010011111001" ,   --120 
    "111110011010010011111001" ,   --121 
    "101001001010010011111001" ,   --122 
    "101100001010010011111001" ,   --123 
    "100110011010010011111001" ,   --124 
    "100100101010010011111001" ,   --125 
    "100000101010010011111001" ,   --126 
    "111110001010010011111001" ,   --127 
    "100000001010010011111001" ,   --128 
    "100100001010010011111001" ,   --129 
    "110000001011000011111001" ,   --130 
    "111110011011000011111001" ,   --131 
    "101001001011000011111001" ,   --132 
    "101100001011000011111001" ,   --133 
    "100110011011000011111001" ,   --134 
    "100100101011000011111001" ,   --135 
    "100000101011000011111001" ,   --136 
    "111110001011000011111001" ,   --137 
    "100000001011000011111001" ,   --138 
    "100100001011000011111001" ,   --139 
    "110000001001100111111001" ,   --140 
    "111110011001100111111001" ,   --141 
    "101001001001100111111001" ,   --142 
    "101100001001100111111001" ,   --143 
    "100110011001100111111001" ,   --144 
    "100100101001100111111001" ,   --145 
    "100000101001100111111001" ,   --146 
    "111110001001100111111001" ,   --147 
    "100000001001100111111001" ,   --148 
    "100100001001100111111001" ,   --149 
    "110000001001001011111001" ,   --150 
    "111110011001001011111001" ,   --151 
    "101001001001001011111001" ,   --152 
    "101100001001001011111001" ,   --153 
    "100110011001001011111001" ,   --154 
    "100100101001001011111001" ,   --155 
    "100000101001001011111001" ,   --156 
    "111110001001001011111001" ,   --157 
    "100000001001001011111001" ,   --158 
    "100100001001001011111001" ,   --159 
    "110000001000001011111001" ,   --160 
    "111110011000001011111001" ,   --161 
    "101001001000001011111001" ,   --162 
    "101100001000001011111001" ,   --163 
    "100110011000001011111001" ,   --164 
    "100100101000001011111001" ,   --165 
    "100000101000001011111001" ,   --166 
    "111110001000001011111001" ,   --167 
    "100000001000001011111001" ,   --168 
    "100100001000001011111001" ,   --169 
    "110000001111100011111001" ,   --170 
    "111110011111100011111001" ,   --171 
    "101001001111100011111001" ,   --172 
    "101100001111100011111001" ,   --173 
    "100110011111100011111001" ,   --174 
    "100100101111100011111001" ,   --175 
    "100000101111100011111001" ,   --176 
    "111110001111100011111001" ,   --177 
    "100000001111100011111001" ,   --178 
    "100100001111100011111001" ,   --179 
    "110000001000000011111001" ,   --180 
    "111110011000000011111001" ,   --181 
    "101001001000000011111001" ,   --182 
    "101100001000000011111001" ,   --183 
    "100110011000000011111001" ,   --184 
    "100100101000000011111001" ,   --185 
    "100000101000000011111001" ,   --186 
    "111110001000000011111001" ,   --187 
    "100000001000000011111001" ,   --188 
    "100100001000000011111001" ,   --189 
    "110000001001000011111001" ,   --190 
    "111110011001000011111001" ,   --191 
    "101001001001000011111001" ,   --192 
    "101100001001000011111001" ,   --193 
    "100110011001000011111001" ,   --194 
    "100100101001000011111001" ,   --195 
    "100000101001000011111001" ,   --196 
    "111110001001000011111001" ,   --197 
    "100000001001000011111001" ,   --198 
    "100100001001000011111001" ,   --199 
    "110000001100000010100100" ,   --200 
    "111110011100000010100100" ,   --201 
    "101001001100000010100100" ,   --202 
    "101100001100000010100100" ,   --203 
    "100110011100000010100100" ,   --204 
    "100100101100000010100100" ,   --205 
    "100000101100000010100100" ,   --206 
    "111110001100000010100100" ,   --207 
    "100000001100000010100100" ,   --208 
    "100100001100000010100100" ,   --209 
    "110000001111100110100100" ,   --210 
    "111110011111100110100100" ,   --211 
    "101001001111100110100100" ,   --212 
    "101100001111100110100100" ,   --213 
    "100110011111100110100100" ,   --214 
    "100100101111100110100100" ,   --215 
    "100000101111100110100100" ,   --216 
    "111110001111100110100100" ,   --217 
    "100000001111100110100100" ,   --218 
    "100100001111100110100100" ,   --219 
    "110000001010010010100100" ,   --220 
    "111110011010010010100100" ,   --221 
    "101001001010010010100100" ,   --222 
    "101100001010010010100100" ,   --223 
    "100110011010010010100100" ,   --224 
    "100100101010010010100100" ,   --225 
    "100000101010010010100100" ,   --226 
    "111110001010010010100100" ,   --227 
    "100000001010010010100100" ,   --228 
    "100100001010010010100100" ,   --229 
    "110000001011000010100100" ,   --230 
    "111110011011000010100100" ,   --231 
    "101001001011000010100100" ,   --232 
    "101100001011000010100100" ,   --233 
    "100110011011000010100100" ,   --234 
    "100100101011000010100100" ,   --235 
    "100000101011000010100100" ,   --236 
    "111110001011000010100100" ,   --237 
    "100000001011000010100100" ,   --238 
    "100100001011000010100100" ,   --239 
    "110000001001100110100100" ,   --240 
    "111110011001100110100100" ,   --241 
    "101001001001100110100100" ,   --242 
    "101100001001100110100100" ,   --243 
    "100110011001100110100100" ,   --244 
    "100100101001100110100100" ,   --245 
    "100000101001100110100100" ,   --246 
    "111110001001100110100100" ,   --247 
    "100000001001100110100100" ,   --248 
    "100100001001100110100100" ,   --249 
    "110000001001001010100100" ,   --250 
    "111110011001001010100100" ,   --251 
    "101001001001001010100100" ,   --252 
    "101100001001001010100100" ,   --253 
    "100110011001001010100100" ,   --254 
    "100100101001001010100100"    --255  
 

  );

begin

  Cur_D_Val_SS_out <= ROM_Data (Cur_D_Val_Out);

end struct;